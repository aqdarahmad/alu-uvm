
include "uvm_macros.svh"
include "sequence_item.sv"
import uvm_pkg::*;
class sequencer extends uvm_Sequencer #(sequence_item);

`uvm_component_utils(sequencer)

// define constructor 
function new(string name = "sequencer",uvm_component parent);
super.new(name , parent);
endfunction :new




endclass : sequencer